
module dispinput(z,o);
 input [3:0]z;
	output reg [13:0]o;
 always @(z)
begin
 case(z)
 4'b0000 : o= 14'b11111110000001;
 4'b0001 : o= 14'b11111111001111;
 4'b0010 : o= 14'b11111110010010;
 4'b0011 : o= 14'b11111110000110;
 4'b0100 : o= 14'b11111111001100;
 4'b0101 : o= 14'b11111110100100;
 4'b0110 : o= 14'b11111110100000;
 4'b0111 : o= 14'b11111110001111;
 4'b1000 : o= 14'b11111110000000;
 4'b1001 : o= 14'b11111110000100;
 4'b1010 : o= 14'b10011110000001;
 4'b1010 : o= 14'b10011111001111;
 4'b1100 : o= 14'b10011110010010;
 4'b1101 : o= 14'b10011110000110;
 4'b1110 : o= 14'b10011111001100;
 4'b1111 : o= 14'b10011110100100;
 
 endcase
 end
 endmodule
 


module dispoutput(p,h);
 input [4:0]p;
 output reg[13:0]h;
 always @(p)
 begin
 case(p)
 5'b00000: h= 14'b11111110000001;
 5'b00001: h= 14'b11111111001111;
 5'b00010: h= 14'b11111110010010;
 5'b00011: h= 14'b11111110000110;
 5'b00100: h= 14'b11111111001100;
 5'b00101: h= 14'b11111110100100;
 5'b00110: h= 14'b11111110100000;
 5'b00111: h= 14'b11111110001111;
 5'b01000: h= 14'b11111110000000;
 5'b01001: h= 14'b11111110000100;
 5'b01010: h= 14'b10011110000001;
 5'b01010: h= 14'b10011111001111;
 5'b01100: h= 14'b10011110010010;
 5'b01101: h= 14'b10011110000110;
 5'b01110: h= 14'b10011111001100;
 5'b01111: h= 14'b10011110100100;
 5'b10000: h= 14'b10011110100000;
 5'b10001: h= 14'b10011110001111;
 5'b10010: h= 14'b10011110000000;
 5'b10011: h= 14'b10011110000100;
 5'b10100: h= 14'b00100100000001;
 5'b10101: h= 14'b00100101001111;
 5'b10110: h= 14'b00100100010010;
 5'b10111: h= 14'b00100100000110;
 5'b11000: h= 14'b00100101001100;
 5'b11001: h= 14'b00100100100100;
 5'b11010: h= 14'b00100100100000;
 5'b11011: h= 14'b00100100001111;
 5'b11100: h= 14'b00100100000000;
 5'b11101: h= 14'b00100100000100;
 5'b11110: h= 14'b00001100000001;
 5'b11111: h= 14'b00001101001111;
 endcase
 end
 endmodule

module Lab5(x,y,cin,sum,d,e,f);
input [3:0] x,y;
input cin;
output reg [4:0] sum;
output [13:0]d ,e,f;

always@(*)
begin
sum = x+y+cin;
end

dispinput firstip(x,d);
dispinput secondip(y,e);
dispoutput sumop(sum,f);
endmodule



